-- Generator Control FPGA
-- DO-254 Compliance
